
`include "single_port_ram.v"
`include "linebuf.v"
`include "linebuf_ram_wrap.v"

`include "linebuf_rgboffset_top.v"
