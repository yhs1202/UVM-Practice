package lb_ro_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "lb_ro_define.sv"

  `include "lb_ro_transfer.sv"
  `include "lb_ro_sequencer.sv"
  `include "lb_ro_driver.sv"
  `include "lb_ro_monitor.sv"
  `include "lb_ro_agent.sv"

  `include "lb_ro_seq_item.sv"
  `include "lb_ro_seq_lib.sv"
  `include "lb_ro_vseq_lib.sv"

endpackage

`include "lb_ro_if.sv"
