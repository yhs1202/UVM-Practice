
import uvm_pkg::*;
`include "uvm_macros.svh"

`include "lb_ro_pkg.sv"
import lb_ro_pkg::*;

`include "lb_ro_if.sv"
`include "lb_ro_sb.sv"
`include "lb_ro_env.sv"

`include "vseqr.sv"
`include "tb.sv"

`include "base_vseq_lib.sv"
`include "base_test.sv"

`include "video_test.sv"

`include "top.sv"
