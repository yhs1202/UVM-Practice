// Agent
class spi_agent extends uvm_agent;
    `uvm_component_utils(spi_agent)

    function new(string name = "agt", uvm_component parent);
        super.new(name, parent);
    endfunction

    uvm_sequencer #(spi_seq_item) sqr;
    spi_driver drv;
    spi_monitor mon;

    function void build_phase(uvm_phase phase);
        super.build_phase(phase);
        sqr = uvm_sequencer#(spi_seq_item)::type_id::create("sqr", this);
        drv = spi_driver::type_id::create("drv", this);
        mon = spi_monitor::type_id::create("mon", this);
    endfunction

    function void connect_phase(uvm_phase phase);
        super.connect_phase(phase);
        drv.seq_item_port.connect(sqr.seq_item_export);
    endfunction
endclass
